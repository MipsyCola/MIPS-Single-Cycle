module Clock_Gen(Clock);
output reg Clock;
initial
begin
Clock=0;
end
always
begin
#31.25
Clock=~(Clock);
end
endmodule
